`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.05.2020 16:09:06
// Design Name: 
// Module Name: Priority_encoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Priority_encoder(
    input [24:0] significand,
    input [7:0] exponent_a,
    output reg [24:0] Significand,
    output [7:0] Exponent_sub
    );
    
    reg [4:0] shift;
    
    always@(significand)
    begin
            casex (significand)
                25'b1_1xxx_xxxx_xxxx_xxxx_xxxx_xxxx :	begin
                                                                Significand = significand;
                                                                shift = 5'd0;
                                                        end 
                25'b1_01xx_xxxx_xxxx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 1;
                                                                shift = 5'd1;
                                                        end
                25'b1_001x_xxxx_xxxx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 2;
                                                                shift = 5'd2;
                                                        end
                25'b1_0001_xxxx_xxxx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 3;
                                                                shift = 5'd3;
                                                        end
                25'b1_0000_1xxx_xxxx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 4;
                                                                shift = 5'd4;
                                                        end
                25'b1_0000_01xx_xxxx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 5;
                                                                shift = 5'd5;
                                                        end
                25'b1_0000_001x_xxxx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 6;
                                                                shift = 5'd6;
                                                        end
                25'b1_0000_0001_xxxx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 7;
                                                                shift = 5'd7;
                                                        end
                25'b1_0000_0000_1xxx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 8;
                                                                shift = 5'd8;
                                                        end
                25'b1_0000_0000_01xx_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 9;
                                                                shift = 5'd9;
                                                        end
                25'b1_0000_0000_001x_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 10;
                                                                shift = 5'd10;
                                                        end
                25'b1_0000_0000_0001_xxxx_xxxx_xxxx :   begin
                                                                Significand = significand << 11;
                                                                shift = 5'd11;
                                                        end
                25'b1_0000_0000_0000_1xxx_xxxx_xxxx :   begin
                                                                Significand = significand << 12;
                                                                shift = 5'd12;
                                                        end
                25'b1_0000_0000_0000_01xx_xxxx_xxxx :   begin
                                                                Significand = significand << 13;
                                                                shift = 5'd13;
                                                        end
                25'b1_0000_0000_0000_001x_xxxx_xxxx :   begin
                                                                Significand = significand << 14;
                                                                shift = 5'd14;
                                                        end
                25'b1_0000_0000_0000_0001_xxxx_xxxx :   begin
                                                                Significand = significand << 15;
                                                                shift = 5'd15;
                                                        end
                25'b1_0000_0000_0000_0000_1xxx_xxxx :   begin
                                                                Significand = significand << 16;
                                                                shift = 5'd16;
                                                        end
                25'b1_0000_0000_0000_0000_01xx_xxxx :   begin
                                                                Significand = significand << 17;
                                                                shift = 5'd17;
                                                        end
                25'b1_0000_0000_0000_0000_001x_xxxx :   begin
                                                                Significand = significand << 18;
                                                                shift = 5'd18;
                                                        end
                25'b1_0000_0000_0000_0000_0001_xxxx :   begin
                                                                Significand = significand << 19;
                                                                shift = 5'd19;
                                                        end
                25'b1_0000_0000_0000_0000_0000_1xxx :   begin
                                                                Significand = significand << 20;
                                                                shift = 5'd20;
                                                        end
                25'b1_0000_0000_0000_0000_0000_01xx :   begin
                                                                Significand = significand << 21;
                                                                shift = 5'd21;
                                                        end
                25'b1_0000_0000_0000_0000_0000_001x :   begin
                                                                Significand = significand << 22;
                                                                shift = 5'd22;
                                                        end
                25'b1_0000_0000_0000_0000_0000_0001 :   begin
                                                                Significand = significand << 23;
                                                                shift = 5'd23;
                                                        end
                25'b1_0000_0000_0000_0000_0000_0000 :   begin
                                                                Significand = significand << 24;
                                                                shift = 5'd24;
                                                        end
                default : 	begin
						Significand = (~significand) + 1'b1;
						shift = 8'd0;
					end
			endcase					                                                shift = 5'd1;
    end  
    assign Exponent_sub = exponent_a - shift;                                                                                                         
endmodule
